module entiremap_rom ( input [10:0]	addr,
						output [79:0]	data
					 );

					  logic [79:0] reg_file[130];  //Instatiating our ROM

always_comb


begin 
                                             //The map will be made of 16x16 blocks so when we do the math
															//the 640X480 screen will be composed of 40x30 of these blocks
															//meaning 40 rows (data_width), 30 columns (amount of data_addr)

reg_file[0]=             80'b111111111111111111111111111111111111111111111111111111111111111111111111111111;
reg_file[1]=             80'b100000000000000000000000000000000000000000000000000000000000000000000000001111;
reg_file[2]=             80'b100000000000000000000000000000000000000000000000000000000000000000000000000111;
reg_file[3]=             80'b100111110001111110001111110001111100001100000001111111000000000111111111100011;
reg_file[4]=             80'b100101010001011010001011010001010100001100000000000000000000000000000000000001;
reg_file[5]=             80'b100111110001111110001111110001111100001100000100000000010000010000000000000001;
reg_file[6]=             80'b100000000000000000000000000000000000001100000100001000010000010001000011100001;
reg_file[7]=             80'b100000000000000000000000000000000000001100000100001000010000010001000000000001;
reg_file[8]=             80'b100110000000000000000001111000000000001100000100001000010000010001000000000001;
reg_file[9]=             80'b100110000000000000000001001000000000001100000100001000010000010001000000000001;
reg_file[10]=            80'b100110011111000011110001111000111110001100000100001000010000010001000111100001;
reg_file[11]=            80'b100110010101000010110000000000101010001100000100001000000000000000000000000001;
reg_file[12]=            80'b100110011011000011010000000000110110001100000100001000000000000000000000000001;
reg_file[13]=            80'b100110010101000010110001111000101010001100000100001000000000000000000110011001;
reg_file[14]=            80'b100110011011000011110001101000110110001100000100000000011111111000100110011001;
reg_file[15]=            80'b100110010101000000000001011000101010001100000100001000000000000000100110011001;
reg_file[16]=            80'b100110011011000000000001101000110110001100000100001000000000000010100110011001;
reg_file[17]=            80'b100110011111000000000001111000111110001000000000000000000000000000100000000001;
reg_file[18]=            80'b100110000000001111110000000000000000001000000000000000000000000000100000000001;
reg_file[19]=            80'b100110000000001010110000000000000000001000000111111111111110000000100000000001;
reg_file[20]=            80'b100110011100001101010000011111000110000000000111111111111110000000100000000001;
reg_file[21]=            80'b100000011100001111110000011111000110000000000000000000000000000000000000000001;
reg_file[22]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[23]=            80'b100000000000000000000000000000000000001000011111111111111111111111111111111001;
reg_file[24]=            80'b100111110001111110001111110001111100001000000000000000000000000000000000000001;
reg_file[25]=            80'b100101010001011010001011010001010100001000000000000000000000000000000000000001;
reg_file[26]=            80'b100111110001111110001111110001111100001000011111111111111111111111111111111001;
reg_file[27]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[28]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[29]=            80'b100111111110011110001111111000111111000001111000011111111111111100001111111001;

reg_file[30]=            80'b100111111110011110001111111000111111000001111000011111111111111100001111111001;
reg_file[31]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[32]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[33]=            80'b100111111111111111111111111111111111110000000111111111100000111111111110000001;
reg_file[34]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[35]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[36]=            80'b100100100001000010010010001000100111111000111100000011111111111111111111111001;
reg_file[37]=            80'b100100100001000010010010001000100110011000101100000010000000111100111011111001;
reg_file[38]=            80'b100100100001000010010010001000100101101000110100000010010100000100001000011001;
reg_file[39]=            80'b100100100001000010010010001000100101101000101100000010000000011100001001111001;
reg_file[40]=            80'b100100100001000010010010001000100110011000110100000010111110000100001000011001;
reg_file[41]=            80'b100100100001000010010010001000100101101000101100000010011100111100111001111001;
reg_file[42]=            80'b100100100001000010010010001000100101101000110100110011111111111111111111111001;
reg_file[43]=            80'b100100100001000010010010001000100110011000101100110000000000000000000000000001;
reg_file[44]=            80'b100100100001000010010010001000100101101000110100110000000000000011100000000001;
reg_file[45]=            80'b100100100001000010010010001000100101101000101100110001110001010100010000000001;
reg_file[46]=            80'b100100100001000010010010001000100110011000110100110010001010110100010000000001;
reg_file[47]=            80'b100000100000000010000010000000100101101000101100000010001000010011010000000001;
reg_file[48]=            80'b100000100000000010000010000000100101101000110100110010001000010000010000000001;
reg_file[49]=            80'b100000100000000010000010000000100110011000101100110001110000010000010000000001;
reg_file[50]=            80'b100000100000000010000010000000100101101000110100000000000000000000000000000001;
reg_file[51]=            80'b100000100000000010000010000000100101101000101100000000000011111111100000000001;
reg_file[52]=            80'b100100100001000010010010001000100110011000110100000000000010000000100000000001;
reg_file[53]=            80'b100100100001000010010010001000100101101000101100000000000010100010100000000001;
reg_file[54]=            80'b100100100001000010010010001000100101101000110100000000000010001000100000000001;
reg_file[55]=            80'b100100100001000010010010001000100110011000101100000000000010010100100000000001;
reg_file[56]=            80'b100000000000000000000000000000000111111000111100000000000011111111100000000001;
reg_file[57]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[58]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[59]=            80'b111111111111111111111111111111111111111111111111111111111111111111111111111111;


/////////////////////////////Map 2

reg_file[70]=            80'b111111111111111111111111111111111111111111111111111111111111111111111111111111;
reg_file[71]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[72]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[73]=            80'b100000111111111111111111111111111110000011111111111111111111111111111111100001;
reg_file[74]=            80'b100000100000000000000000000000000000000000000000000000000000000000000000100001;
reg_file[75]=            80'b100000100000000000000000000000000000000000000000000000000000000000000000100001;
reg_file[76]=            80'b100000100000111111111111111111111111111111111111111111111111111111110000100001;
reg_file[77]=            80'b100000100000100000000000000000000000000000000000000000000000000000010000100001; 
reg_file[78]=            80'b100000100000100000000000000000000000000000000000000000000000000000010000100001;
reg_file[79]=            80'b100000100000100011111111111111111110000011111111111111111111111000010000100001;
reg_file[80]=            80'b100000100000100010000000000000000000000000000000000000000000001000010000100001;
reg_file[81]=            80'b100000100000100010000000000000000000000000000000000000000000001000010000100001;
reg_file[82]=            80'b100000100000100010011111111111111111111111111111111111111110001000010000100001;
reg_file[83]=            80'b100000100000000010000000000000000000000000000000000000000000001000010000000001;
reg_file[84]=            80'b100000100000000010000000000000000000000000000000000000000000001000010000000001;
reg_file[85]=            80'b100000100000100010011111111111111110000111111111111111111110001000010000100001;
reg_file[86]=            80'b100000100000100010000000000000000000000000000000000000000000001000010000100001;
reg_file[87]=            80'b100000100000100010000000000000000000000000000000000000000000001000010000100001;
reg_file[88]=            80'b100000100000100011111111111111111111111111111111111111111111111000010000100001;
reg_file[89]=            80'b100000100000100000000000000000000000000000000000000000000000000000010000100001;
reg_file[90]=            80'b100000100000100000000000000000000000000000000000000000000000000000010000100001;
reg_file[91]=            80'b100000100000111111111111111111111110000111111111111111111111111111110000100001;
reg_file[92]=            80'b100000100000000000000000000000000000000000000000000000000000000000000000100001;
reg_file[93]=            80'b100000100000000000000000000000000000000000000000000000000000000000000000100001;
reg_file[94]=            80'b100000100000000000000000000000000000000000000000000000000000000000000000100001;
reg_file[95]=            80'b100000111111111111111111111111111111111111111111111111111111111111111111100001;
reg_file[96]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[97]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[98]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[99]=            80'b100111111110011110001111111000111111000001111000011111111111111100001111111001;

reg_file[100]=            80'b100111111110011110001111111000111111000001111000011111111111111100001111111001;
reg_file[101]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[102]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[103]=            80'b100111111111111111111111111111111111110000000111111111100000111111111110000001;
reg_file[104]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[105]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[106]=            80'b100100100001000010010010001000100111111000111111111111111111111111111111111001;
reg_file[107]=            80'b100100100001000010010010001000100110011000101100000010000000111100111011111001;
reg_file[108]=            80'b100100100001000010010010001000100101101000110100000010010100000100001000011001;
reg_file[109]=            80'b100100100001000010010010001000100101101000101100000010000000011100001001111001;
reg_file[110]=            80'b100100100001000010010010001000100110011000110100110010111110000100001000011001;
reg_file[111]=            80'b100100100001000010010010001000100101101000101100110010011100111100111001111001;
reg_file[112]=            80'b100100100001000010010010001000100101101000110100110011111111111111111111111001;
reg_file[113]=            80'b100100100001000010010010001000100110011000101100110000000000000000000000000001;
reg_file[114]=            80'b100100100001000010010010001000100000000000110100110000000000000000000000000001;
reg_file[115]=            80'b100100100001000010010010001000100000000000101100110000000000000000000000000001;
reg_file[116]=            80'b100100100001000010010010001000011111111111111100110000000000000000000000000001;
reg_file[117]=            80'b100100100000000010000010000000000000000000000000110000000000000000000000010001;
reg_file[118]=            80'b100100100000000010000010000000000000000000000000110000000000000000000000010001;
reg_file[119]=            80'b100100100000000010000010000000000000000000000000110000000000000000000000010001;
reg_file[120]=            80'b100100100000000010000010000000111111111111111100110000000000000000000000010001;
reg_file[121]=            80'b100100000000000010000010000000100000000000101100110001111111111111111111110001;
reg_file[122]=            80'b100100000001000000010000001000100000000000110100110001100110000000100000010001;
reg_file[123]=            80'b100100000001000000010000001000100111111000101100000001011010100010101001010001;
reg_file[124]=            80'b100100000001000000010000001000100101101000110100000001011010001000110000110001;
reg_file[125]=            80'b100111111111111111111111111111100110011000101100000001100110010100100110010001;
reg_file[126]=            80'b100000000000000000000000000000000111111000111111111111111111111111111111110001;
reg_file[127]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[128]=            80'b100000000000000000000000000000000000000000000000000000000000000000000000000001;
reg_file[129]=            80'b111111111111111111111111111111111111111111111111111111111111111111111111111111;


end

assign data = reg_file[addr];



endmodule 